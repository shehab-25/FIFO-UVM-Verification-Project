package shared_pkg;
    parameter FIFO_WIDTH = 16;
    parameter FIFO_DEPTH = 8;
    int RD_EN_ON_DIST = 50;
    int WR_EN_ON_DIST = 50;
endpackage